module IF_stage#
(
    parameter handler_addr = 32'd1000
)
(
    ID_PFC, EX_PFC, PC_src, inst_mem_in, PC_write, clk, inst, rst
);
	
input [31:0] ID_PFC, EX_PFC;
input [2:0] PC_src;
input PC_write, clk, rst;

output [31:0] inst;
inout [31:0] inst_mem_in;

wire [31:0] pc_reg_in;


MUX_8x1 PC_src_mux(inst_mem_in + 1'b1, handler_addr, ID_PFC, inst_mem_in, EX_PFC, 0, 0, 0, PC_src, pc_reg_in);

PC_register pc_reg(pc_reg_in, inst_mem_in, PC_write, clk, rst); 

IM inst_mem(inst_mem_in , inst, clk);

endmodule

module RS();



endmodule



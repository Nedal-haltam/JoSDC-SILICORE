
module control_unit(opcode, regwrite, memread, memwrite);

   input [6:0] 	opcode;
	
	output reg			regwrite; 																
	output reg			memread; 								
	output reg			memwrite;
	
	
parameter add = 7'h20, sub = 7'h22, addu = 7'h21, subu = 7'h23, addi = 7'h48, and_ = 7'h24, andi = 7'h4c, or_ = 7'h25, ori = 7'h4d, xor_ = 7'h26, 
		    xori = 7'h4e, nor_ = 7'h27, sll = 7'h00, srl = 7'h02, lw = 7'h63, sw = 7'h6b, beq = 7'h44, bne = 7'h45, blt = 7'h50, bge = 7'h51, 
			 j = 7'h42, jal = 7'h43, jr = 7'h08, slt = 7'h2a, hlt_inst = 7'b1111111;

	
	
always @(opcode) begin
		{regwrite, memread, memwrite} <= 0; //By Default all Control Signals are equal to zero
		// if none of these instructions then the the regwrite = 1
		if (!(opcode == jr || opcode == sw || opcode == beq || opcode == bne || opcode == blt || opcode == bge || opcode == j))
			regwrite <= 1'b1;
		if (opcode == lw)
			memread <= 1'b1;
		if (opcode == sw)
			memwrite <= 1'b1;
			
end	
endmodule




module OOO_CPU
(
    input input_clk, rst,
    output reg [31:0] cycles_consumed
);

`include "opcodes.txt"

wire [31:0] PC, PC_out, Branch_Target_Addr;
wire PC_src, clk;
// InstQ
wire [ 11:0] InstQ_opcode;
wire [3:0] InstQ_ALUOP;
wire [ 4:0] InstQ_rs, InstQ_rt, InstQ_rd, InstQ_shamt;
wire [15:0] InstQ_immediate;
wire [25:0] InstQ_address;
wire InstQ_VALID_Inst;


// RegFile
wire [31:0] RegFile_RP1_Reg1, RegFile_RP1_Reg2;
wire [4:0] RegFile_RP1_Reg1_ROBEN, RegFile_RP1_Reg2_ROBEN;


// ROB
wire ROB_FULL_FLAG;
wire ROB_EXCEPTION_Flag;
wire ROB_FLUSH_Flag;
wire [11:0] ROB_Commit_opcode;
wire [4:0] ROB_Commit_Rd;
wire [31:0] ROB_Commit_Write_Data;
wire [2:0] ROB_Commit_Control_Signals;
wire [4:0] ROB_Start_Index;
wire [4:0] ROB_End_Index;
wire [31:0] ROB_RP1_Write_Data1, ROB_RP1_Write_Data2;
wire ROB_RP1_Ready1, ROB_RP1_Ready2;


// RS
wire RS_FULL_FLAG;
wire [4:0] RS_FU_RS_ID, RS_FU_ROBEN;
wire [11:0] RS_FU_opcode;
wire [3:0] RS_FU_ALUOP;
wire [31:0] RS_FU_Val1, RS_FU_Val2;
wire [31:0] RS_FU_Immediate;


// FU
wire [31:0] FU_Result;
wire [4:0] FU_ROBEN;
wire [11:0] FU_opcode;
wire FU_Is_Free;



// Address Unit
wire AU_LdStB_VALID_Inst;
wire [4:0]  AU_LdStB_ROBEN;
wire [4:0]  AU_LdStB_Rd;
wire [11:0] AU_LdStB_opcode;
wire [4:0]  AU_LdStB_ROBEN1, AU_LdStB_ROBEN2;
wire [31:0] AU_LdStB_ROBEN1_VAL, AU_LdStB_ROBEN2_VAL;
wire [31:0] AU_LdStB_Immediate;
wire [31:0] AU_LdStB_EA, AU_LdStB_Write_Data;


// Load Store Buffer
wire LdStB_MEMU_VALID_Inst;
wire [4:0]  LdStB_MEMU_ROBEN;
wire [4:0]  LdStB_MEMU_Rd;
wire [11:0] LdStB_MEMU_opcode;
wire [4:0]  LdStB_MEMU_ROBEN1, LdStB_MEMU_ROBEN2;
wire [31:0] LdStB_MEMU_ROBEN1_VAL, LdStB_MEMU_ROBEN2_VAL;
wire [31:0] LdStB_MEMU_Immediate;
wire [31:0] LdStB_MEMU_EA, LdStB_MEMU_Write_Data;
wire [3:0] LdStB_Start_Index;
wire [3:0] LdStB_End_Index;

// Memory Unit
wire [4:0] MEMU_ROBEN;
wire [31:0] MEMU_Result;



// CDB
wire [4:0] CDB_ROBEN1;
wire [31:0] CDB_Write_Data1;
wire [4:0] CDB_ROBEN2;
wire [31:0] CDB_Write_Data2;






wire hlt;
assign hlt = ROB_Commit_opcode == hlt_inst;
nor hlt_logic(clk, input_clk, hlt);


always@(negedge clk , posedge rst) begin
	if (rst)
		cycles_consumed <= 32'd0;
	else
		cycles_consumed <= cycles_consumed + 32'd1;
end


/*
PC_src_mux:
    - change the PC_src value based on decoded or commit instruction
TODO:
    - consider: j, jal, jr
    - what about FULL ROB what will happen
*/
assign PC = (ROB_FLUSH_Flag == 1'b1) ? ROB_Commit_Write_Data :
(
    (InstQ_opcode == hlt_inst) ? PC_out : 
    (
        (InstQ_opcode == beq || InstQ_opcode == bne) ? PC_out + {{16{InstQ_immediate[15]}},InstQ_immediate} : PC_out + 1'b1
    )
);
// assign PC = (PC_src) ? Branch_Target_Addr : PC_out + 1'b1;


PC_register pcreg(PC, PC_out, ~ROB_FULL_FLAG || ROB_FLUSH_Flag , clk, rst);

InstQ instq
(
    .clk(clk), 
    .rst(rst),
    .PC(PC_out),
    
    .opcode(InstQ_opcode),
    .rs(InstQ_rs), 
    .rt(InstQ_rt), 
    .rd(InstQ_rd), 
    .shamt(InstQ_shamt),
    .immediate(InstQ_immediate),
    .address(InstQ_address),
    .VALID_Inst(InstQ_VALID_Inst)
);

reg ROB_HLT;
always@(posedge clk, posedge rst) begin
    if (rst)
        ROB_HLT = 1'b1;
    else
        ROB_HLT = InstQ_opcode == hlt_inst;
end

RegFile regfile
(
    .clk(clk),
    .rst(rst),

    .WP1_Wen(ROB_Commit_Control_Signals[2]), 
    .Decoded_WP1_Wen((!(InstQ_opcode == jr || InstQ_opcode == sw || InstQ_opcode == beq || 
                        InstQ_opcode == bne || InstQ_opcode == j))),
    .WP1_ROBEN
    (
        (ROB_Start_Index == 5'd1) ? 5'd16 : (ROB_Start_Index - 1'b1)
    ), 
    .Decoded_WP1_ROBEN
    (
        (ROB_FULL_FLAG || ROB_FLUSH_Flag) ? 5'd0 : ROB_End_Index
    ), 
    .WP1_DRindex(ROB_Commit_Rd), 
    .Decoded_WP1_DRindex
    (
        (InstQ_opcode == jal) ? 5'd31 : 
        (
            (InstQ_opcode[11:6] == 6'd0) ? InstQ_rd : InstQ_rt
        )
    ), 
    .WP1_Data(ROB_Commit_Write_Data),

    // inputs
    .RP1_index1(InstQ_rs), 
    .RP1_index2(InstQ_rt),
    // outputs
    .RP1_Reg1(RegFile_RP1_Reg1), 
    .RP1_Reg2(RegFile_RP1_Reg2),
    .RP1_Reg1_ROBEN(RegFile_RP1_Reg1_ROBEN), 
    .RP1_Reg2_ROBEN(RegFile_RP1_Reg2_ROBEN)
);



ROB rob
(
    .clk(clk), 
    .rst(rst),
    .Decoded_opcode(InstQ_opcode),
    .Decoded_Rd
    (
        (InstQ_opcode == addi || InstQ_opcode == andi || InstQ_opcode == ori || InstQ_opcode == xori || 
         InstQ_opcode == sll  || InstQ_opcode == srl  || InstQ_opcode == slti || InstQ_opcode == lw) ? InstQ_rt : InstQ_rd
    ),
    .Decoded_prediction(InstQ_opcode == beq | InstQ_opcode == bne),
    .Branch_Target_Addr(PC_out + 1'b1),

    // TODO: get the rest of the sources
    .CDB_ROBEN1(CDB_ROBEN1),
    .CDB_ROBEN1_Write_Data(CDB_Write_Data1),

    .CDB_ROBEN2(CDB_ROBEN2),
    .CDB_ROBEN2_Write_Data(CDB_Write_Data2),
    .CDB_Branch_Decision(FU_Branch_Decision),

    .VALID_Inst
    (
        ~rst && ~ROB_HLT && ~ROB_FLUSH_Flag && ~ROB_FULL_FLAG 
    ),

    .FULL_FLAG(ROB_FULL_FLAG),
    .EXCEPTION_Flag(ROB_EXCEPTION_Flag),
    .FLUSH_Flag(ROB_FLUSH_Flag),

    .Commit_opcode(ROB_Commit_opcode),
    .Commit_Rd(ROB_Commit_Rd),
    .Commit_Write_Data(ROB_Commit_Write_Data),
    .Commit_Control_Signals(ROB_Commit_Control_Signals),

    .RP1_ROBEN1(RegFile_RP1_Reg1_ROBEN), 
    .RP1_ROBEN2(RegFile_RP1_Reg2_ROBEN),

    .RP1_Write_Data1(ROB_RP1_Write_Data1), 
    .RP1_Write_Data2(ROB_RP1_Write_Data2),
    .RP1_Ready1(ROB_RP1_Ready1), 
    .RP1_Ready2(ROB_RP1_Ready2),

    .Start_Index(ROB_Start_Index),
    .End_Index(ROB_End_Index)
);


ALU_OPER alu_op(InstQ_opcode, InstQ_ALUOP);

RS rs
(
    .clk(clk), 
    .rst(rst),
    .opcode(InstQ_opcode),
    .ALUOP(InstQ_ALUOP),
    .ROBEN((ROB_End_Index == 5'd1) ? 5'd16 : (ROB_End_Index - 1'b1)),
    .ROBEN1
    (
        (RegFile_RP1_Reg1_ROBEN == 0) ? 5'd0 : 
        (
            (ROB_RP1_Ready1) ? 5'd0 : RegFile_RP1_Reg1_ROBEN
        )
    ), 
    .ROBEN2
    (
        (InstQ_opcode == addi || InstQ_opcode == andi || InstQ_opcode == ori || InstQ_opcode == xori || 
         InstQ_opcode == sll  || InstQ_opcode == srl  || InstQ_opcode == slti) ? 5'd0 : 
         (
            (RegFile_RP1_Reg2_ROBEN == 0) ? 5'd0 : 
            (
                (ROB_RP1_Ready2) ? 5'd0 : RegFile_RP1_Reg2_ROBEN
            )
         )
    ), 
    .ROBEN1_VAL
    (
        (RegFile_RP1_Reg1_ROBEN == 0) ? RegFile_RP1_Reg1 : ROB_RP1_Write_Data1
    ), 
    .ROBEN2_VAL
    (
        (RegFile_RP1_Reg2_ROBEN == 0) ? RegFile_RP1_Reg2 : ROB_RP1_Write_Data2
    ), 
    .Immediate
    (
        (InstQ_opcode == sll || InstQ_opcode == srl) ? {27'd0,InstQ_shamt} : 
        (
            (InstQ_opcode == andi || InstQ_opcode == ori || InstQ_opcode == xori) ? {16'd0,InstQ_immediate} : 
            (
                {{16{InstQ_immediate[15]}},InstQ_immediate}
            )
        )
    ),
    // TODO: get the rest of the sources
    .CDB_ROBEN1(CDB_ROBEN1),
    .CDB_ROBEN1_VAL(CDB_Write_Data1),
    .CDB_ROBEN2(CDB_ROBEN2),
    .CDB_ROBEN2_VAL(CDB_Write_Data2),

    .VALID_Inst
    (
        InstQ_opcode != hlt_inst && InstQ_VALID_Inst && ~ROB_FULL_FLAG && ~ROB_FLUSH_Flag && InstQ_opcode != lw && InstQ_opcode != sw
    ),
    .FU_Is_Free(FU_Is_Free),

    .FULL_FLAG(RS_FULL_FLAG),

    .RS_FU_RS_ID(RS_FU_RS_ID),
    .RS_FU_ROBEN(RS_FU_ROBEN),
    .RS_FU_opcode(RS_FU_opcode),   
    .RS_FU_ALUOP(RS_FU_ALUOP),
    .RS_FU_Val1(RS_FU_Val1), 
    .RS_FU_Val2(RS_FU_Val2),
    .RS_FU_Immediate(RS_FU_Immediate)

);

ALU alu
(
    .clk(clk),
    .rst(rst),
    .ROBEN(RS_FU_ROBEN),
    .opcode(RS_FU_opcode),
    .A(RS_FU_Val1), 
    .B
    (
        (RS_FU_opcode == addi || RS_FU_opcode == andi || RS_FU_opcode == ori || RS_FU_opcode == xori || 
         RS_FU_opcode == sll  || RS_FU_opcode == srl  || RS_FU_opcode == slti) ? RS_FU_Immediate : RS_FU_Val2
    ), 
    .ALUOP(RS_FU_ALUOP),

    .FU_res(FU_Result), 
    .FU_Branch_Decision(FU_Branch_Decision),
    .FU_ROBEN(FU_ROBEN),
    .FU_opcode(FU_opcode),
    .FU_Is_Free(FU_Is_Free)
);




CDB cdb
(
    .ROBEN1(FU_ROBEN),
    .Write_Data1(FU_Result),

    .ROBEN2(MEMU_ROBEN),
    .Write_Data2(MEMU_Result),

    // input [4:0] ROBEN3,
    // input [31:0] Write_Data3,

    // input [4:0] ROBEN4,
    // input [31:0] Write_Data4,


    .out_ROBEN1(CDB_ROBEN1),
    .out_Write_Data1(CDB_Write_Data1),

    .out_ROBEN2(CDB_ROBEN2),
    .out_Write_Data2(CDB_Write_Data2)

    // output [4:0] out_ROBEN3,
    // output [31:0] out_Write_Data3,

    // output [4:0] out_ROBEN4,
    // output [31:0] out_Write_Data4
);



AddressUnit AU
(
    .Decoded_ROBEN(ROB_End_Index - 1'b1),
    .Decoded_Rd(InstQ_rt),
    .Decoded_opcode(InstQ_opcode),
    .ROBEN1
    (
        (RegFile_RP1_Reg1_ROBEN == 0) ? 5'd0 : 
        (
            (ROB_RP1_Ready1) ? 5'd0 : RegFile_RP1_Reg1_ROBEN
        )
    ), 
    .ROBEN2
    (
        (InstQ_opcode == lw) ? 5'd0 : 
        (
            (RegFile_RP1_Reg2_ROBEN == 0) ? 5'd0 : 
            (
                (ROB_RP1_Ready2) ? 5'd0 : RegFile_RP1_Reg2_ROBEN
            )
        )
    ),
    .ROBEN1_VAL
    (
        (RegFile_RP1_Reg1_ROBEN == 0) ? RegFile_RP1_Reg1 : ROB_RP1_Write_Data1
    ), 
    .ROBEN2_VAL
    (
        (RegFile_RP1_Reg2_ROBEN == 0) ? RegFile_RP1_Reg2 : ROB_RP1_Write_Data2
    ), 
    .Immediate({{16{InstQ_immediate[15]}},InstQ_immediate}),


    .AU_LdStB_VALID_Inst(AU_LdStB_VALID_Inst),
    .AU_LdStB_ROBEN(AU_LdStB_ROBEN),
    .AU_LdStB_Rd(AU_LdStB_Rd),
    .AU_LdStB_opcode(AU_LdStB_opcode),
    .AU_LdStB_ROBEN1(AU_LdStB_ROBEN1), 
    .AU_LdStB_ROBEN2(AU_LdStB_ROBEN2),
    .AU_LdStB_ROBEN1_VAL(AU_LdStB_ROBEN1_VAL), 
    .AU_LdStB_ROBEN2_VAL(AU_LdStB_ROBEN2_VAL),
    .AU_LdStB_Immediate(AU_LdStB_Immediate),
    .AU_LdStB_EA(AU_LdStB_EA)
);



/*
TOOD: 
    - we may separate the LdSt Buffer to load buffer and store buffer but two things should be taken into consideration
        
        - for both lw, sw we should forward the needed registers (lw: register to calc EA, sw: register to calc EA, and another to store in the MEM)
        so if the register is available there is no problem otherwise:
            - case 1: we take the ROBEN from the ROB
        
        - secondly: (lw,sw) memory dependencies through similar EA 
        we should check for similar EA once we enter the load/store buffers if we are `ready`
        or once the needed register for calc the EA is forwarded to us from the CDB.
        we should find the last sw that wants to write on the same EA 
        and based on him we take its register and call ourself `ready` or take its ROBEN if its unavailable and wait for it
            we care about the following three cases if there is similar EAs
            - RAW: we forward the register to be written to the memory from the store instruction or take its ROBEN.......
            - WAW:
            - WAR:
*/
LdStBuffer ldstbuffer
(
    .clk(clk), 
    .rst(rst),
    .VALID_Inst(AU_LdStB_VALID_Inst),
    .ROBEN(AU_LdStB_ROBEN),
    .Rd(AU_LdStB_Rd),
    .opcode(AU_LdStB_opcode),
    .ROBEN1(AU_LdStB_ROBEN1), 
    .ROBEN2(AU_LdStB_ROBEN2),
    .ROBEN1_VAL(AU_LdStB_ROBEN1_VAL), 
    .ROBEN2_VAL(AU_LdStB_ROBEN2_VAL),
    .Immediate(AU_LdStB_Immediate),
    .EA(AU_LdStB_EA),

    .CDB_ROBEN(CDB_ROBEN1),
    .CDB_ROBEN_VAL(CDB_Write_Data1),


    .out_VALID_Inst(LdStB_MEMU_VALID_Inst),
    .out_ROBEN(LdStB_MEMU_ROBEN),
    .out_Rd(LdStB_MEMU_Rd),
    .out_opcode(LdStB_MEMU_opcode),
    .out_ROBEN1(LdStB_MEMU_ROBEN1), 
    .out_ROBEN2(LdStB_MEMU_ROBEN2),
    .out_ROBEN1_VAL(LdStB_MEMU_ROBEN1_VAL), 
    .out_ROBEN2_VAL(LdStB_MEMU_ROBEN2_VAL),
    .out_Immediate(LdStB_MEMU_Immediate),
    .out_EA(LdStB_MEMU_EA),

    .Start_Index(LdStB_Start_Index),
    .End_Index(LdStB_End_Index)
);


DM datamemory
(
    .clk(clk), 
    .ROBEN((LdStB_MEMU_VALID_Inst) ? LdStB_MEMU_ROBEN : 5'd0),
    .Read_en
    (
        (LdStB_MEMU_VALID_Inst) ? LdStB_MEMU_opcode == lw : 1'b0
    ), 
    .Write_en
    (
        (LdStB_MEMU_VALID_Inst) ? LdStB_MEMU_opcode == sw : 1'b0
    ), 
    .address(LdStB_MEMU_EA),
    .data(LdStB_MEMU_ROBEN2_VAL),

    .MEMU_ROBEN(MEMU_ROBEN),
    .MEMU_Result(MEMU_Result)

);



/*
TODO:
    - MemoryUnit
    - CDB
*/






endmodule
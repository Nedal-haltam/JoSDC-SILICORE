module BranchController();


// output PCsrc;

endmodule
 





module RS();



endmodule



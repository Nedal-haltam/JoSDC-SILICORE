module InstQ
(
    input clk, rst,
    input  [31:0] PC,
    
    output reg [ 11:0] opcode,
    output reg [ 4:0] rs, rt, rd, shamt,
    output reg [15:0] immediate,
    output reg [25:0] address,
    output reg VALID_Inst
);


reg [31:0] InstMem [63:0];

wire [31:0] inst;

assign inst = InstMem[PC];


always@(negedge clk, posedge rst) begin
    if (rst) begin
        opcode <= 0;
        rs <= 0;
        rt <= 0;
        rd <= 0;
        shamt <= 0;
        immediate <= 0;
        address <= 0;
        VALID_Inst <= 1'b0;
    end
    else begin
        if (inst[31:26] == 0)
            opcode    <= { inst[31:26], inst[5:0] };
        else
            opcode    <= { inst[31:26], 6'd0 };

        rs        <= inst[25:21];
        rt        <= inst[20:16];
        rd        <= inst[15:11];
        shamt     <= inst[10:6];
        immediate <= inst[15:0];
        address   <= inst[25:0];
        VALID_Inst <= 1'b1;
    end
end



initial begin


InstMem[  0] <= 32'h200100FF; // addi $1 $zero 255
InstMem[  1] <= 32'h20420001; // addi $2 $2 1
InstMem[  2] <= 32'h00000000; // nop
InstMem[  3] <= 32'h1441FFFE; // bne $2 $1 -2
InstMem[  4] <= 32'hFC000000; // hlt




// InstMem[  0] <= 32'h20010064; // addi $1 $zero 100
// InstMem[  1] <= 32'h2042000A; // addi $2 $2 10
// InstMem[  2] <= 32'h10220002; // beq $1 $2 2
// InstMem[  3] <= 32'h1042FFFE; // beq $2 $2 -2
// InstMem[  4] <= 32'hFC000000; // hlt






/* run the following to simulate in VS Code, note you should be in '\GitHub Repos\JoSDC-SILICORE\SSOOO' in the terminal
> iverilog -o sim -D vscode .\OOO_CPU_Sim.v
> vvp sim
*/







end


endmodule


`include "RS.v"

module RS_tb();



endmodule



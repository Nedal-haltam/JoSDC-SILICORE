
`define HALF_CYCLE 1
`define ONE_CLK (2 * `HALF_CYCLE)
`define ADVANCE_N_CYCLE(N) #(`ONE_CLK * N);

`define MAX_CLOCKS (100 * 1000 * 1000)
`define reset 2 * `ONE_CLK


`ifndef vscode
`timescale 1ns/1ps
`endif


`define MEMORY_SIZE 2048
`define MEMORY_BITS 11
`define ROB_SIZE_bits (4)
`define BUFFER_SIZE_bitslsbuffer (4)
`define BUFFER_SIZE_bitsRS (4)
`define ROB_SIZE ((1 << `ROB_SIZE_bits))

`ifdef vscode

`include "./AddressUnit&ld_st buffer/AddressUnit.v"
`include "./AddressUnit&ld_st buffer/LSBuffer.v"
`include "./Common Data Bus/CDB.v"
`include "./Instruction Queue/InstQ.v"
`include "./Memory Unit/DM.v"
`include "./Register File/RegFile.v"
`include "./Reorder Buffer/ROB.v"
`include "./Reservation Station/RS.v"
`include "./Functional Unit/compare_equal.v"
`include "./Functional Unit/ALU_OPER.v"
`include "./Functional Unit/ALU.v"
`include "PC_register.v"
`include "BranchPredictor.v"
`include "SSOOO_CPU.v"

`endif

module SSOOO_Sim();

reg clk = 0, rst = 0;
wire [31 : 0] cycles_consumed, StallCount;
`ifdef vscode
wire real BranchPredictionCount, BranchPredictionMissCount;
`else
wire [31:0] BranchPredictionCount, BranchPredictionMissCount;
`endif

SSOOO_CPU #(.CORE_SELECT(1'b0)) cpu
(
	.input_clk(clk), 
	.rst(rst),
    .cycles_consumed(cycles_consumed),
    .StallCount(StallCount),
    .BranchPredictionCount(BranchPredictionCount),
    .BranchPredictionMissCount(BranchPredictionMissCount)
);


always #(`HALF_CYCLE) clk <= ~clk;
initial begin

`ifdef VCD_OUT

$dumpfile(`VCD_OUT);
$dumpvars;

`else

// $dumpfile("SSOOO_Waveform.vcd");
// $dumpvars;

`endif

rst <= 1; #(`reset) rst <= 0;

#(`MAX_CLOCKS + 1);
$display("\t\tNumber of cycles consumed: %d", cycles_consumed);
$display("\t\tStallCount: %d", StallCount);
$display("\t\tExecuted Instruction   Count: %d", cycles_consumed - StallCount);
$display("\t\tBranch Prediction      Count: %d", BranchPredictionCount);
$display("\t\tBranch Prediction HIT  Count: %d", BranchPredictionCount - BranchPredictionMissCount);
$display("\t\tBranch Prediction HIT  Rate : %.3f%%", ((BranchPredictionCount - BranchPredictionMissCount) / BranchPredictionCount) * 100);
$display("\t\tBranch Prediction Miss Count: %d", BranchPredictionMissCount);
$display("\t\tBranch Prediction Miss Rate : %.3f%%", (BranchPredictionMissCount / BranchPredictionCount) * 100);



$finish;

end

endmodule


/*


//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module SSOOO_CPU(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW
);



//=======================================================
//  REG/WIRE declarations
//=======================================================




//=======================================================
//  Structural coding
//=======================================================



endmodule
*/
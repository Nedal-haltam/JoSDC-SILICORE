module DM(addr , Data_In , Data_Out , WR , clk);

parameter bit_width = 32;
input [bit_width - 1:0] addr , Data_In;
input WR , clk;
output [bit_width - 1:0] Data_Out;

reg [bit_width - 1:0] data_mem [255 : 0];
  
always@ (posedge clk)  
  if (WR == 1'b1)
    data_mem[addr] = Data_In;

assign Data_Out = data_mem[addr];




`ifdef sim
initial begin
  #(`timeunits + `reset);
  // iterating through some of the addresses of the memory to check if the program loaded and stored the values properly
  $display("Reading Data Memory Content : ");
  for (integer i = 50; i >= 0; i = i - 1)
    $display("addr = %d , Mem[addr] = %d",i,$signed(data_mem[i]));

end 
`endif
      
endmodule
module MUX_F_8();




endmodule